** Profile: "SCHEMATIC1-trnasiente"  [ C:\Users\Leonan\Google Drive\UFRJ\Projeto Final\simulacoes\Orcad\instrumentacao\instrumentacao-pspicefiles\schematic1\trnasiente.sim ] 

** Creating circuit file "trnasiente.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 1u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
